module Register32(
	in,
	out,
	clk,
	en
);

endmodule