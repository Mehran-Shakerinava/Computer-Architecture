module SingleCycleCPU;


Register32 PC(
	
);



endmodule