module Adder(
	a,
	b,
	out
);


endmodule