module RAM(
	write_addr,
	read_addr,
	en,
	write_data,
	read_data,
	clk
);

endmodule